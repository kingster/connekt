[ambari-server]
10.33.109.42

[ac]
10.33.253.88
10.33.157.7
10.34.93.241
10.33.121.23
10.32.153.197
10.33.25.217
10.33.105.242
10.32.45.230
10.34.1.246
10.32.169.215
10.32.1.231
10.32.133.186
10.32.33.222
10.32.73.234
10.32.85.23
10.32.17.229
10.32.65.239
10.32.61.232
10.34.97.18
